    Mac OS X            	   2  �     �                                    ATTR     �   �   �                  �     com.apple.lastuseddate#PS       �   �  "com.apple.LaunchServices.OpenWith    o��e    C@�    bplist00�WversionTpath_bundleidentifier _!/System/Applications/TextEdit.app_com.apple.TextEdit/1U                            j                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              This resource fork intentionally left blank                                                                                                                                                                                                                            ��